##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Wed Jun  8 12:06:42 2022
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 1900.720000 BY 2339.200000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 115.825 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 618.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1105 LAYER met4  ;
    ANTENNAMAXAREACAR 10.1559 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 51.6564 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.154225 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 5.050000 0.000000 5.350000 0.800000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 89.7106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 478.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 80.5261 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1.550000 0.000000 1.850000 0.800000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.550000 0.000000 396.850000 0.800000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.150000 0.000000 133.450000 0.800000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.350000 0.000000 400.650000 0.800000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 392.650000 0.000000 392.950000 0.800000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 388.850000 0.000000 389.150000 0.800000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 385.050000 0.000000 385.350000 0.800000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 381.250000 0.000000 381.550000 0.800000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 255.350000 0.000000 255.650000 0.800000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 251.450000 0.000000 251.750000 0.800000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 247.750000 0.000000 248.050000 0.800000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 243.850000 0.000000 244.150000 0.800000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 240.150000 0.000000 240.450000 0.800000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.250000 0.000000 236.550000 0.800000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.350000 0.000000 232.650000 0.800000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 228.650000 0.000000 228.950000 0.800000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 224.850000 0.000000 225.150000 0.800000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.950000 0.000000 221.250000 0.800000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.150000 0.000000 217.450000 0.800000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.350000 0.000000 213.650000 0.800000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.550000 0.000000 209.850000 0.800000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.750000 0.000000 206.050000 0.800000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850000 0.000000 202.150000 0.800000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 198.150000 0.000000 198.450000 0.800000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.250000 0.000000 194.550000 0.800000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 190.550000 0.000000 190.850000 0.800000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.650000 0.000000 186.950000 0.800000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.750000 0.000000 183.050000 0.800000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 179.050000 0.000000 179.350000 0.800000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 175.250000 0.000000 175.550000 0.800000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 171.350000 0.000000 171.650000 0.800000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 167.550000 0.000000 167.850000 0.800000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 163.750000 0.000000 164.050000 0.800000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 160.050000 0.000000 160.350000 0.800000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.150000 0.000000 156.450000 0.800000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.250000 0.000000 152.550000 0.800000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.550000 0.000000 148.850000 0.800000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.750000 0.000000 145.050000 0.800000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.850000 0.000000 141.150000 0.800000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 137.050000 0.000000 137.350000 0.800000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.450000 0.000000 129.750000 0.800000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.650000 0.000000 125.950000 0.800000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.750000 0.000000 122.050000 0.800000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.950000 0.000000 118.250000 0.800000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 114.150000 0.000000 114.450000 0.800000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.450000 0.000000 110.750000 0.800000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.550000 0.000000 106.850000 0.800000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.650000 0.000000 102.950000 0.800000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 98.950000 0.000000 99.250000 0.800000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.150000 0.000000 95.450000 0.800000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.250000 0.000000 91.550000 0.800000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.450000 0.000000 87.750000 0.800000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.550000 0.000000 83.850000 0.800000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.950000 0.000000 80.250000 0.800000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.050000 0.000000 76.350000 0.800000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.150000 0.000000 72.450000 0.800000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.350000 0.000000 68.650000 0.800000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.650000 0.000000 64.950000 0.800000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.750000 0.000000 61.050000 0.800000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.950000 0.000000 57.250000 0.800000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.050000 0.000000 53.350000 0.800000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.350000 0.000000 49.650000 0.800000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.550000 0.000000 45.850000 0.800000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.650000 0.000000 41.950000 0.800000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 37.850000 0.000000 38.150000 0.800000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 34.050000 0.000000 34.350000 0.800000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.250000 0.000000 30.550000 0.800000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.450000 0.000000 26.750000 0.800000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.550000 0.000000 22.850000 0.800000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.750000 0.000000 19.050000 0.800000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 15.050000 0.000000 15.350000 0.800000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 11.150000 0.000000 11.450000 0.800000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 7.350000 0.000000 7.650000 0.800000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 377.450000 0.000000 377.750000 0.800000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 373.550000 0.000000 373.850000 0.800000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 369.750000 0.000000 370.050000 0.800000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 365.950000 0.000000 366.250000 0.800000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 362.150000 0.000000 362.450000 0.800000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 358.350000 0.000000 358.650000 0.800000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 354.450000 0.000000 354.750000 0.800000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 350.750000 0.000000 351.050000 0.800000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 346.950000 0.000000 347.250000 0.800000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 343.050000 0.000000 343.350000 0.800000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 339.250000 0.000000 339.550000 0.800000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 335.450000 0.000000 335.750000 0.800000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 331.550000 0.000000 331.850000 0.800000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 327.850000 0.000000 328.150000 0.800000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 323.950000 0.000000 324.250000 0.800000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 320.250000 0.000000 320.550000 0.800000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 316.350000 0.000000 316.650000 0.800000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 312.550000 0.000000 312.850000 0.800000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 308.750000 0.000000 309.050000 0.800000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 304.950000 0.000000 305.250000 0.800000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 301.150000 0.000000 301.450000 0.800000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 297.350000 0.000000 297.650000 0.800000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 293.450000 0.000000 293.750000 0.800000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 289.650000 0.000000 289.950000 0.800000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 285.850000 0.000000 286.150000 0.800000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 281.950000 0.000000 282.250000 0.800000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 278.250000 0.000000 278.550000 0.800000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 274.350000 0.000000 274.650000 0.800000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 270.650000 0.000000 270.950000 0.800000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 266.750000 0.000000 267.050000 0.800000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 262.950000 0.000000 263.250000 0.800000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.377 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 621.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 259.150000 0.000000 259.450000 0.800000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 888.650000 0.000000 888.950000 0.800000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 884.750000 0.000000 885.050000 0.800000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 880.950000 0.000000 881.250000 0.800000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 877.150000 0.000000 877.450000 0.800000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 873.450000 0.000000 873.750000 0.800000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 869.550000 0.000000 869.850000 0.800000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 865.650000 0.000000 865.950000 0.800000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 861.950000 0.000000 862.250000 0.800000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.150000 0.000000 858.450000 0.800000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 854.250000 0.000000 854.550000 0.800000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 850.450000 0.000000 850.750000 0.800000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.650000 0.000000 846.950000 0.800000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 842.850000 0.000000 843.150000 0.800000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 839.050000 0.000000 839.350000 0.800000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.150000 0.000000 835.450000 0.800000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 831.450000 0.000000 831.750000 0.800000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 827.550000 0.000000 827.850000 0.800000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 823.750000 0.000000 824.050000 0.800000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.950000 0.000000 820.250000 0.800000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 816.150000 0.000000 816.450000 0.800000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 812.350000 0.000000 812.650000 0.800000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 808.550000 0.000000 808.850000 0.800000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 804.650000 0.000000 804.950000 0.800000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 800.850000 0.000000 801.150000 0.800000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 797.050000 0.000000 797.350000 0.800000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 793.250000 0.000000 793.550000 0.800000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 789.450000 0.000000 789.750000 0.800000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 785.550000 0.000000 785.850000 0.800000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 781.850000 0.000000 782.150000 0.800000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 777.950000 0.000000 778.250000 0.800000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 774.150000 0.000000 774.450000 0.800000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 770.350000 0.000000 770.650000 0.800000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 766.550000 0.000000 766.850000 0.800000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 762.750000 0.000000 763.050000 0.800000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 758.950000 0.000000 759.250000 0.800000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 755.050000 0.000000 755.350000 0.800000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 751.350000 0.000000 751.650000 0.800000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 747.450000 0.000000 747.750000 0.800000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 743.650000 0.000000 743.950000 0.800000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 739.850000 0.000000 740.150000 0.800000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 736.050000 0.000000 736.350000 0.800000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 732.250000 0.000000 732.550000 0.800000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 728.350000 0.000000 728.650000 0.800000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 724.550000 0.000000 724.850000 0.800000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 720.750000 0.000000 721.050000 0.800000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 716.950000 0.000000 717.250000 0.800000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 713.050000 0.000000 713.350000 0.800000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 709.350000 0.000000 709.650000 0.800000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 705.450000 0.000000 705.750000 0.800000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 701.750000 0.000000 702.050000 0.800000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 697.850000 0.000000 698.150000 0.800000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 694.050000 0.000000 694.350000 0.800000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 690.250000 0.000000 690.550000 0.800000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 686.450000 0.000000 686.750000 0.800000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 682.650000 0.000000 682.950000 0.800000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 678.750000 0.000000 679.050000 0.800000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.950000 0.000000 675.250000 0.800000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 671.250000 0.000000 671.550000 0.800000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 667.350000 0.000000 667.650000 0.800000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 663.450000 0.000000 663.750000 0.800000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 659.750000 0.000000 660.050000 0.800000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 655.950000 0.000000 656.250000 0.800000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 652.150000 0.000000 652.450000 0.800000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 648.250000 0.000000 648.550000 0.800000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 644.450000 0.000000 644.750000 0.800000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 640.650000 0.000000 640.950000 0.800000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 636.850000 0.000000 637.150000 0.800000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 632.950000 0.000000 633.250000 0.800000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 629.150000 0.000000 629.450000 0.800000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 625.350000 0.000000 625.650000 0.800000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 621.650000 0.000000 621.950000 0.800000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 617.750000 0.000000 618.050000 0.800000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.850000 0.000000 614.150000 0.800000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 610.150000 0.000000 610.450000 0.800000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 606.350000 0.000000 606.650000 0.800000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 602.450000 0.000000 602.750000 0.800000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 598.650000 0.000000 598.950000 0.800000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 594.850000 0.000000 595.150000 0.800000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 591.150000 0.000000 591.450000 0.800000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.250000 0.000000 587.550000 0.800000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350000 0.000000 583.650000 0.800000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 579.550000 0.000000 579.850000 0.800000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 575.850000 0.000000 576.150000 0.800000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 572.050000 0.000000 572.350000 0.800000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 568.150000 0.000000 568.450000 0.800000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 564.250000 0.000000 564.550000 0.800000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 560.550000 0.000000 560.850000 0.800000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 556.750000 0.000000 557.050000 0.800000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 552.850000 0.000000 553.150000 0.800000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 549.050000 0.000000 549.350000 0.800000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 545.250000 0.000000 545.550000 0.800000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 541.550000 0.000000 541.850000 0.800000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 537.650000 0.000000 537.950000 0.800000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 533.750000 0.000000 534.050000 0.800000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 529.950000 0.000000 530.250000 0.800000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 526.250000 0.000000 526.550000 0.800000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 522.350000 0.000000 522.650000 0.800000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 518.550000 0.000000 518.850000 0.800000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 514.650000 0.000000 514.950000 0.800000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 511.050000 0.000000 511.350000 0.800000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 507.150000 0.000000 507.450000 0.800000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 503.250000 0.000000 503.550000 0.800000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 499.450000 0.000000 499.750000 0.800000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 495.750000 0.000000 496.050000 0.800000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 491.950000 0.000000 492.250000 0.800000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 488.050000 0.000000 488.350000 0.800000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 484.150000 0.000000 484.450000 0.800000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 480.450000 0.000000 480.750000 0.800000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.650000 0.000000 476.950000 0.800000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 472.750000 0.000000 473.050000 0.800000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 468.950000 0.000000 469.250000 0.800000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 465.150000 0.000000 465.450000 0.800000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 8.91071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.1525 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 461.450000 0.000000 461.750000 0.800000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 8.90687 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.5626 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 457.550000 0.000000 457.850000 0.800000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 6.23913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.5429 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.335662 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 453.650000 0.000000 453.950000 0.800000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 11.4418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.8657 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.24303 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 449.850000 0.000000 450.150000 0.800000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 9.44713 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.3545 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 446.150000 0.000000 446.450000 0.800000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 9.24424 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.3323 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 442.250000 0.000000 442.550000 0.800000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 8.18631 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.8494 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 438.450000 0.000000 438.750000 0.800000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 9.43879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.1586 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 434.550000 0.000000 434.850000 0.800000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 6.17174 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 27.6583 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 430.850000 0.000000 431.150000 0.800000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 10.1741 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.8636 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 427.050000 0.000000 427.350000 0.800000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 6.84322 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.2831 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.311653 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 423.150000 0.000000 423.450000 0.800000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 9.19333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.0778 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 419.350000 0.000000 419.650000 0.800000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 8.01688 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.0248 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 415.550000 0.000000 415.850000 0.800000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 9.57919 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.5101 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 411.750000 0.000000 412.050000 0.800000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.55616 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.8626 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.261549 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 407.950000 0.000000 408.250000 0.800000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 10.82 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.1943 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.330009 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 404.050000 0.000000 404.350000 0.800000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.66 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.1 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1376.850000 0.000000 1377.150000 0.800000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1373.150000 0.000000 1373.450000 0.800000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.66 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.1 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1369.350000 0.000000 1369.650000 0.800000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1365.450000 0.000000 1365.750000 0.800000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1361.650000 0.000000 1361.950000 0.800000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1357.850000 0.000000 1358.150000 0.800000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1354.150000 0.000000 1354.450000 0.800000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1350.250000 0.000000 1350.550000 0.800000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1346.350000 0.000000 1346.650000 0.800000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1342.650000 0.000000 1342.950000 0.800000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1338.750000 0.000000 1339.050000 0.800000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1335.050000 0.000000 1335.350000 0.800000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1331.150000 0.000000 1331.450000 0.800000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1327.350000 0.000000 1327.650000 0.800000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1323.550000 0.000000 1323.850000 0.800000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1319.750000 0.000000 1320.050000 0.800000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1315.850000 0.000000 1316.150000 0.800000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1312.050000 0.000000 1312.350000 0.800000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1308.250000 0.000000 1308.550000 0.800000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1304.550000 0.000000 1304.850000 0.800000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1300.650000 0.000000 1300.950000 0.800000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1296.750000 0.000000 1297.050000 0.800000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1293.050000 0.000000 1293.350000 0.800000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1289.150000 0.000000 1289.450000 0.800000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1285.350000 0.000000 1285.650000 0.800000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1281.550000 0.000000 1281.850000 0.800000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1277.750000 0.000000 1278.050000 0.800000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1273.950000 0.000000 1274.250000 0.800000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1270.150000 0.000000 1270.450000 0.800000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1266.250000 0.000000 1266.550000 0.800000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1262.550000 0.000000 1262.850000 0.800000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1258.650000 0.000000 1258.950000 0.800000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1254.950000 0.000000 1255.250000 0.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1251.050000 0.000000 1251.350000 0.800000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1247.250000 0.000000 1247.550000 0.800000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1243.450000 0.000000 1243.750000 0.800000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1239.550000 0.000000 1239.850000 0.800000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1235.750000 0.000000 1236.050000 0.800000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1231.950000 0.000000 1232.250000 0.800000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1228.150000 0.000000 1228.450000 0.800000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1224.350000 0.000000 1224.650000 0.800000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1220.550000 0.000000 1220.850000 0.800000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1216.650000 0.000000 1216.950000 0.800000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1212.950000 0.000000 1213.250000 0.800000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1209.050000 0.000000 1209.350000 0.800000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1205.250000 0.000000 1205.550000 0.800000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1201.450000 0.000000 1201.750000 0.800000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1197.650000 0.000000 1197.950000 0.800000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1193.850000 0.000000 1194.150000 0.800000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1189.950000 0.000000 1190.250000 0.800000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1186.150000 0.000000 1186.450000 0.800000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1182.450000 0.000000 1182.750000 0.800000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1178.550000 0.000000 1178.850000 0.800000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.595 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1174.650000 0.000000 1174.950000 0.800000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1170.950000 0.000000 1171.250000 0.800000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1167.150000 0.000000 1167.450000 0.800000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1163.350000 0.000000 1163.650000 0.800000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1159.450000 0.000000 1159.750000 0.800000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1155.650000 0.000000 1155.950000 0.800000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1151.850000 0.000000 1152.150000 0.800000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1148.050000 0.000000 1148.350000 0.800000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1144.250000 0.000000 1144.550000 0.800000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1140.350000 0.000000 1140.650000 0.800000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1136.550000 0.000000 1136.850000 0.800000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1132.850000 0.000000 1133.150000 0.800000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1128.950000 0.000000 1129.250000 0.800000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1125.050000 0.000000 1125.350000 0.800000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1121.350000 0.000000 1121.650000 0.800000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1117.550000 0.000000 1117.850000 0.800000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1113.750000 0.000000 1114.050000 0.800000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1109.850000 0.000000 1110.150000 0.800000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1106.050000 0.000000 1106.350000 0.800000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1102.350000 0.000000 1102.650000 0.800000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1098.450000 0.000000 1098.750000 0.800000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1094.550000 0.000000 1094.850000 0.800000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1090.750000 0.000000 1091.050000 0.800000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1087.050000 0.000000 1087.350000 0.800000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1083.250000 0.000000 1083.550000 0.800000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1079.350000 0.000000 1079.650000 0.800000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1075.450000 0.000000 1075.750000 0.800000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1071.750000 0.000000 1072.050000 0.800000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1067.950000 0.000000 1068.250000 0.800000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1064.150000 0.000000 1064.450000 0.800000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1060.250000 0.000000 1060.550000 0.800000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1056.450000 0.000000 1056.750000 0.800000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1052.750000 0.000000 1053.050000 0.800000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1048.850000 0.000000 1049.150000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1044.950000 0.000000 1045.250000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1041.150000 0.000000 1041.450000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1037.450000 0.000000 1037.750000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1033.650000 0.000000 1033.950000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1029.750000 0.000000 1030.050000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1025.850000 0.000000 1026.150000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1022.250000 0.000000 1022.550000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1018.350000 0.000000 1018.650000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1014.450000 0.000000 1014.750000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1010.650000 0.000000 1010.950000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1006.950000 0.000000 1007.250000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1003.150000 0.000000 1003.450000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 999.250000 0.000000 999.550000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 995.350000 0.000000 995.650000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 991.650000 0.000000 991.950000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 987.850000 0.000000 988.150000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 983.950000 0.000000 984.250000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 980.150000 0.000000 980.450000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 976.350000 0.000000 976.650000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 972.650000 0.000000 972.950000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 968.750000 0.000000 969.050000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 964.850000 0.000000 965.150000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 961.050000 0.000000 961.350000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 957.350000 0.000000 957.650000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 953.550000 0.000000 953.850000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 949.650000 0.000000 949.950000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 945.750000 0.000000 946.050000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 942.050000 0.000000 942.350000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 938.250000 0.000000 938.550000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 934.350000 0.000000 934.650000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 930.550000 0.000000 930.850000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 926.750000 0.000000 927.050000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 923.050000 0.000000 923.350000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 919.150000 0.000000 919.450000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 915.250000 0.000000 915.550000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 911.550000 0.000000 911.850000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 907.750000 0.000000 908.050000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 903.850000 0.000000 904.150000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 900.050000 0.000000 900.350000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.8474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 896.250000 0.000000 896.550000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.7574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 505.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 892.450000 0.000000 892.750000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1865.350000 0.000000 1865.650000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1861.450000 0.000000 1861.750000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1857.550000 0.000000 1857.850000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1853.850000 0.000000 1854.150000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1850.050000 0.000000 1850.350000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1846.250000 0.000000 1846.550000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1842.350000 0.000000 1842.650000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1838.550000 0.000000 1838.850000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1834.750000 0.000000 1835.050000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1830.950000 0.000000 1831.250000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1827.150000 0.000000 1827.450000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1823.250000 0.000000 1823.550000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1819.450000 0.000000 1819.750000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1815.750000 0.000000 1816.050000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1811.850000 0.000000 1812.150000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1807.950000 0.000000 1808.250000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1804.250000 0.000000 1804.550000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1800.450000 0.000000 1800.750000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.650000 0.000000 1796.950000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1792.750000 0.000000 1793.050000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1788.950000 0.000000 1789.250000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1785.150000 0.000000 1785.450000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.350000 0.000000 1781.650000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1777.450000 0.000000 1777.750000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1773.750000 0.000000 1774.050000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1769.850000 0.000000 1770.150000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1766.150000 0.000000 1766.450000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1762.250000 0.000000 1762.550000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1758.450000 0.000000 1758.750000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1754.650000 0.000000 1754.950000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1750.850000 0.000000 1751.150000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1746.950000 0.000000 1747.250000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1743.150000 0.000000 1743.450000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1739.350000 0.000000 1739.650000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1735.550000 0.000000 1735.850000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1731.750000 0.000000 1732.050000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1727.850000 0.000000 1728.150000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1724.150000 0.000000 1724.450000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1720.250000 0.000000 1720.550000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1716.550000 0.000000 1716.850000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1712.650000 0.000000 1712.950000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1708.850000 0.000000 1709.150000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1705.050000 0.000000 1705.350000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1701.250000 0.000000 1701.550000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1697.350000 0.000000 1697.650000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1693.650000 0.000000 1693.950000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1689.750000 0.000000 1690.050000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1685.950000 0.000000 1686.250000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1682.150000 0.000000 1682.450000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1678.350000 0.000000 1678.650000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1674.550000 0.000000 1674.850000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1670.650000 0.000000 1670.950000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1666.850000 0.000000 1667.150000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1663.050000 0.000000 1663.350000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1659.250000 0.000000 1659.550000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1655.450000 0.000000 1655.750000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1651.650000 0.000000 1651.950000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1647.750000 0.000000 1648.050000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1644.050000 0.000000 1644.350000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1640.150000 0.000000 1640.450000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1636.350000 0.000000 1636.650000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1632.550000 0.000000 1632.850000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1628.750000 0.000000 1629.050000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1624.950000 0.000000 1625.250000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1621.050000 0.000000 1621.350000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1617.250000 0.000000 1617.550000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1613.550000 0.000000 1613.850000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1609.650000 0.000000 1609.950000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1605.850000 0.000000 1606.150000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1602.050000 0.000000 1602.350000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1598.250000 0.000000 1598.550000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1594.450000 0.000000 1594.750000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1590.550000 0.000000 1590.850000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1586.650000 0.000000 1586.950000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1582.950000 0.000000 1583.250000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1579.150000 0.000000 1579.450000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1575.350000 0.000000 1575.650000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1571.450000 0.000000 1571.750000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1567.650000 0.000000 1567.950000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1563.950000 0.000000 1564.250000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1560.050000 0.000000 1560.350000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1556.150000 0.000000 1556.450000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1552.450000 0.000000 1552.750000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1548.650000 0.000000 1548.950000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1544.850000 0.000000 1545.150000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1540.950000 0.000000 1541.250000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1537.050000 0.000000 1537.350000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1533.450000 0.000000 1533.750000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1529.550000 0.000000 1529.850000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1525.750000 0.000000 1526.050000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1521.850000 0.000000 1522.150000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1518.150000 0.000000 1518.450000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1514.350000 0.000000 1514.650000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1510.450000 0.000000 1510.750000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1506.550000 0.000000 1506.850000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1502.850000 0.000000 1503.150000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1499.050000 0.000000 1499.350000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1495.250000 0.000000 1495.550000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1491.350000 0.000000 1491.650000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1487.550000 0.000000 1487.850000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1483.850000 0.000000 1484.150000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1479.950000 0.000000 1480.250000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1476.050000 0.000000 1476.350000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1472.250000 0.000000 1472.550000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1468.550000 0.000000 1468.850000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1464.750000 0.000000 1465.050000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1460.850000 0.000000 1461.150000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1456.950000 0.000000 1457.250000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1453.350000 0.000000 1453.650000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1449.450000 0.000000 1449.750000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1445.650000 0.000000 1445.950000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1441.750000 0.000000 1442.050000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1437.950000 0.000000 1438.250000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1434.250000 0.000000 1434.550000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1430.350000 0.000000 1430.650000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1426.450000 0.000000 1426.750000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1422.750000 0.000000 1423.050000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1418.950000 0.000000 1419.250000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1415.150000 0.000000 1415.450000 0.800000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1411.250000 0.000000 1411.550000 0.800000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1407.450000 0.000000 1407.750000 0.800000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1403.750000 0.000000 1404.050000 0.800000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1399.850000 0.000000 1400.150000 0.800000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1395.950000 0.000000 1396.250000 0.800000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1392.150000 0.000000 1392.450000 0.800000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1388.350000 0.000000 1388.650000 0.800000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1384.650000 0.000000 1384.950000 0.800000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1380.750000 0.000000 1381.050000 0.800000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8259 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 70.7349 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.889 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 87.015000 0.800000 87.415000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5574 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 9.76455 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 51.0094 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 217.840000 0.800000 218.240000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3514 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.164 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 348.940000 0.800000 349.340000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4525 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 62.7024 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 331.706 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 523.465000 0.800000 523.865000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.521 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 215.702 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1141.01 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.27222 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 698.080000 0.800000 698.480000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9555 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 10.6932 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 62.7793 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 872.605000 0.800000 873.005000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.737 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 19.4843 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 109.826 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1047.220000 0.800000 1047.620000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3939 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 16.927 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 76.2381 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1221.835000 0.800000 1222.235000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 29.3984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.111 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1396.360000 0.800000 1396.760000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7875 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 59.154 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.762 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1570.975000 0.800000 1571.375000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.227 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 20.3716 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.878 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1745.590000 0.800000 1745.990000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1920.210000 0.800000 1920.610000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.845 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 26.5476 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.079 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2094.730000 0.800000 2095.130000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6384 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 91.1587 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2269.440000 0.800000 2269.840000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.1936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.6264 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 100.053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.905 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 107.250000 2338.400000 107.550000 2339.200000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 70.3143 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 343.214 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 322.150000 2338.400000 322.450000 2339.200000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4663 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2183 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.397 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 537.150000 2338.400000 537.450000 2339.200000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 124.165 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 637.817 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 752.250000 2338.400000 752.550000 2339.200000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 49.2706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 967.250000 2338.400000 967.550000 2339.200000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 98.7071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.659 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1182.150000 2338.400000 1182.450000 2339.200000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 117.187 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 585.119 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1397.150000 2338.400000 1397.450000 2339.200000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1832 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 51.173 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.779 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1612.150000 2338.400000 1612.450000 2339.200000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 39.6056 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 188.5 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1827.150000 2338.400000 1827.450000 2339.200000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.623 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 542.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 579.051 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3065.99 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2224.085000 1900.720000 2224.485000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.5953 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 335.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 518.667 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2762.99 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2046.155000 1900.720000 2046.555000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.792 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5119 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.127 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1868.230000 1900.720000 1868.630000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 61.6415 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1690.210000 1900.720000 1690.610000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.3852 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 149.831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 708.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1512.280000 1900.720000 1512.680000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 42.9341 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 211.063 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1334.350000 1900.720000 1334.750000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 56.7397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.087 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1156.330000 1900.720000 1156.730000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9479 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 138.949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 719.892 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 978.405000 1900.720000 978.805000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 800.475000 1900.720000 800.875000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1289 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 154.248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 798.468 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 666.985000 1900.720000 667.385000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 533.585000 1900.720000 533.985000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.804 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 389.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 610.842 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3245.17 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 400.090000 1900.720000 400.490000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2814 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 19.6929 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.7698 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 266.600000 1900.720000 267.000000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.7224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 157.994 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 753.921 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 133.110000 1900.720000 133.510000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 10.840000 1900.720000 11.240000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.5647 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 382.624 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 43.315000 0.800000 43.715000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 156.245 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 835.192 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 174.325000 0.800000 174.725000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 107.417 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 574.776 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 305.240000 0.800000 305.640000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 109.218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 583.44 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 479.855000 0.800000 480.255000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.3622 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 493.544 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 654.380000 0.800000 654.780000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 171.235 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 916.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 308.27 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1644.46 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854141 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 828.995000 0.800000 829.395000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.9944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 347.112 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1003.610000 0.800000 1004.010000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.6586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 416.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 334.575 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1791.54 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.94505 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1178.230000 0.800000 1178.630000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1352.845000 0.800000 1353.245000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.3722 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.264 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1527.460000 0.800000 1527.860000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.2057 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 423.376 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1702.075000 0.800000 1702.475000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.896 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1876.600000 0.800000 1877.000000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 140.122 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 748.736 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2051.215000 0.800000 2051.615000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 246.49 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1315.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 671.464 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3571.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2225.830000 0.800000 2226.230000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 217.547 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1160.72 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 53.450000 2338.400000 53.750000 2339.200000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 268.450000 2338.400000 268.750000 2339.200000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8181 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 LAYER met3  ;
    ANTENNAMAXAREACAR 100.956 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 520.108 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.790972 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 483.450000 2338.400000 483.750000 2339.200000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 698.450000 2338.400000 698.750000 2339.200000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 93.4774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 499.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.9687 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 272.98 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1456.83 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3915 LAYER met4  ;
    ANTENNAMAXAREACAR 754.342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3982.51 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.46806 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 913.350000 2338.400000 913.650000 2339.200000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 149.552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 797.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.534 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 261.245 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1393.78 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3915 LAYER met4  ;
    ANTENNAMAXAREACAR 733.252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3882.9 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.873787 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1128.450000 2338.400000 1128.750000 2339.200000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1343.450000 2338.400000 1343.750000 2339.200000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1558.450000 2338.400000 1558.750000 2339.200000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1773.350000 2338.400000 1773.650000 2339.200000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.2784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.96 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2268.610000 1900.720000 2269.010000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.1502 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 375.08 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2090.590000 1900.720000 2090.990000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0989 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.336 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1912.665000 1900.720000 1913.065000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.24 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1734.830000 1900.720000 1735.230000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.7994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.072 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1556.810000 1900.720000 1557.210000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.1842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.928 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1378.790000 1900.720000 1379.190000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.904 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1200.770000 1900.720000 1201.170000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 129.078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 690.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8215 LAYER met4  ;
    ANTENNAMAXAREACAR 158.83 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 803.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.485815 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1022.930000 1900.720000 1023.330000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3215 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.984 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 845.005000 1900.720000 845.405000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 129.018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 689.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8215 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7266 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.418 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 711.510000 1900.720000 711.910000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.3344 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.112 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 578.020000 1900.720000 578.420000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.9472 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 432.664 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 444.530000 1900.720000 444.930000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.349 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 504.344 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 311.130000 1900.720000 311.530000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.3849 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.528 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 177.545000 1900.720000 177.945000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.349 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 504.344 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 44.235000 1900.720000 44.635000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 154.585 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 825.4 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 4.030000 0.800000 4.430000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 298.51 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1593.47 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 130.625000 0.800000 131.025000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 239.532 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1278.92 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 261.630000 0.800000 262.030000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 645.04 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 436.155000 0.800000 436.555000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.1192 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 428.248 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 610.770000 0.800000 611.170000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.9732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 454.136 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 785.390000 0.800000 785.790000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.4702 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.12 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 960.005000 0.800000 960.405000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.1194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.112 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1134.530000 0.800000 1134.930000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.6667 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.168 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1309.145000 0.800000 1309.545000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.696 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1483.760000 0.800000 1484.160000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.6887 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.952 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1658.375000 0.800000 1658.775000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.216 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1832.900000 0.800000 1833.300000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8297 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.704 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2007.515000 0.800000 2007.915000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8979 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.264 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2182.225000 0.800000 2182.625000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 5.850000 2338.400000 6.150000 2339.200000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.1454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 214.750000 2338.400000 215.050000 2339.200000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 429.650000 2338.400000 429.950000 2339.200000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 644.650000 2338.400000 644.950000 2339.200000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.5392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 350.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 859.650000 2338.400000 859.950000 2339.200000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 108.925 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 581.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1074.650000 2338.400000 1074.950000 2339.200000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1289.550000 2338.400000 1289.850000 2339.200000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1504.650000 2338.400000 1504.950000 2339.200000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1719.650000 2338.400000 1719.950000 2339.200000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2849 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.328 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2307.345000 1900.720000 2307.745000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0912 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.432 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2135.120000 1900.720000 2135.520000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6626 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.872 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1957.100000 1900.720000 1957.500000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6199 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.448 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1779.265000 1900.720000 1779.665000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.0699 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.848 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1601.245000 1900.720000 1601.645000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7199 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.648 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1423.315000 1900.720000 1423.715000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2512 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.952 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1245.390000 1900.720000 1245.790000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.261 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 546.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4095 LAYER met4  ;
    ANTENNAMAXAREACAR 275.233 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1457.67 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.397379 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1067.370000 1900.720000 1067.770000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 129.078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 690.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8215 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7479 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.701 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 889.440000 1900.720000 889.840000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.33 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 546.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4095 LAYER met4  ;
    ANTENNAMAXAREACAR 249.889 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1334.39 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 756.040000 1900.720000 756.440000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 129.078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 690.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8215 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7479 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.701 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 622.550000 1900.720000 622.950000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.1049 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.368 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 489.055000 1900.720000 489.455000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 143.628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 766.696 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 355.565000 1900.720000 355.965000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.2814 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.976 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 222.070000 1900.720000 222.470000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 143.628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 766.696 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 88.670000 1900.720000 89.070000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 392.455000 0.800000 392.855000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 567.070000 0.800000 567.470000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 741.690000 0.800000 742.090000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 916.210000 0.800000 916.610000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1090.920000 0.800000 1091.320000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1265.535000 0.800000 1265.935000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1440.150000 0.800000 1440.550000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1614.675000 0.800000 1615.075000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1789.290000 0.800000 1789.690000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 1963.910000 0.800000 1964.310000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2138.525000 0.800000 2138.925000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2306.425000 0.800000 2306.825000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 160.950000 2338.400000 161.250000 2339.200000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.050000 2338.400000 376.350000 2339.200000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.950000 2338.400000 591.250000 2339.200000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 805.950000 2338.400000 806.250000 2339.200000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1020.850000 2338.400000 1021.150000 2339.200000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1235.950000 2338.400000 1236.250000 2339.200000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1450.850000 2338.400000 1451.150000 2339.200000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1665.850000 2338.400000 1666.150000 2339.200000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1873.650000 2338.400000 1873.950000 2339.200000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2179.555000 1900.720000 2179.955000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 2001.630000 1900.720000 2002.030000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1823.700000 1900.720000 1824.100000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1645.770000 1900.720000 1646.170000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1467.750000 1900.720000 1468.150000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1289.825000 1900.720000 1290.225000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 1111.805000 1900.720000 1112.205000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1899.920000 933.970000 1900.720000 934.370000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1869.050000 0.000000 1869.350000 0.800000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1878.250000 0.000000 1878.550000 0.800000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.64 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1875.550000 0.000000 1875.850000 0.800000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 225.692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1204.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.464 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1872.850000 0.000000 1873.150000 0.800000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1888.480000 8.060000 1892.480000 2330.460000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.780000 8.060000 11.780000 2330.460000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1191.640000 1860.520000 1193.380000 2255.300000 ;
      LAYER met3 ;
        RECT 716.320000 1860.520000 1193.380000 1862.260000 ;
      LAYER met3 ;
        RECT 716.320000 2253.560000 1193.380000 2255.300000 ;
      LAYER met4 ;
        RECT 716.320000 1860.520000 718.060000 2255.300000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1191.640000 1363.020000 1193.380000 1757.800000 ;
      LAYER met3 ;
        RECT 716.320000 1363.020000 1193.380000 1364.760000 ;
      LAYER met3 ;
        RECT 716.320000 1756.060000 1193.380000 1757.800000 ;
      LAYER met4 ;
        RECT 716.320000 1363.020000 718.060000 1757.800000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1191.640000 865.520000 1193.380000 1260.300000 ;
      LAYER met3 ;
        RECT 716.320000 865.520000 1193.380000 867.260000 ;
      LAYER met3 ;
        RECT 716.320000 1258.560000 1193.380000 1260.300000 ;
      LAYER met4 ;
        RECT 716.320000 865.520000 718.060000 1260.300000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1191.640000 368.020000 1193.380000 762.800000 ;
      LAYER met3 ;
        RECT 716.320000 368.020000 1193.380000 369.760000 ;
      LAYER met3 ;
        RECT 716.320000 761.060000 1193.380000 762.800000 ;
      LAYER met4 ;
        RECT 716.320000 368.020000 718.060000 762.800000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1821.420000 1860.520000 1823.160000 2255.300000 ;
      LAYER met3 ;
        RECT 1346.100000 1860.520000 1823.160000 1862.260000 ;
      LAYER met3 ;
        RECT 1346.100000 2253.560000 1823.160000 2255.300000 ;
      LAYER met4 ;
        RECT 1346.100000 1860.520000 1347.840000 2255.300000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1821.420000 1363.020000 1823.160000 1757.800000 ;
      LAYER met3 ;
        RECT 1346.100000 1363.020000 1823.160000 1364.760000 ;
      LAYER met3 ;
        RECT 1346.100000 1756.060000 1823.160000 1757.800000 ;
      LAYER met4 ;
        RECT 1346.100000 1363.020000 1347.840000 1757.800000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1821.420000 865.520000 1823.160000 1260.300000 ;
      LAYER met3 ;
        RECT 1346.100000 865.520000 1823.160000 867.260000 ;
      LAYER met3 ;
        RECT 1346.100000 1258.560000 1823.160000 1260.300000 ;
      LAYER met4 ;
        RECT 1346.100000 865.520000 1347.840000 1260.300000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1821.420000 368.020000 1823.160000 762.800000 ;
      LAYER met3 ;
        RECT 1346.100000 368.020000 1823.160000 369.760000 ;
      LAYER met3 ;
        RECT 1346.100000 761.060000 1823.160000 762.800000 ;
      LAYER met4 ;
        RECT 1346.100000 368.020000 1347.840000 762.800000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1882.480000 14.060000 1886.480000 2324.460000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.780000 14.060000 17.780000 2324.460000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 719.720000 2250.160000 1189.980000 2251.900000 ;
      LAYER met3 ;
        RECT 719.720000 1863.920000 1189.980000 1865.660000 ;
      LAYER met4 ;
        RECT 719.720000 1863.920000 721.460000 2251.900000 ;
      LAYER met4 ;
        RECT 1188.240000 1863.920000 1189.980000 2251.900000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 719.720000 1752.660000 1189.980000 1754.400000 ;
      LAYER met3 ;
        RECT 719.720000 1366.420000 1189.980000 1368.160000 ;
      LAYER met4 ;
        RECT 719.720000 1366.420000 721.460000 1754.400000 ;
      LAYER met4 ;
        RECT 1188.240000 1366.420000 1189.980000 1754.400000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 719.720000 1255.160000 1189.980000 1256.900000 ;
      LAYER met3 ;
        RECT 719.720000 868.920000 1189.980000 870.660000 ;
      LAYER met4 ;
        RECT 719.720000 868.920000 721.460000 1256.900000 ;
      LAYER met4 ;
        RECT 1188.240000 868.920000 1189.980000 1256.900000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 719.720000 757.660000 1189.980000 759.400000 ;
      LAYER met3 ;
        RECT 719.720000 371.420000 1189.980000 373.160000 ;
      LAYER met4 ;
        RECT 719.720000 371.420000 721.460000 759.400000 ;
      LAYER met4 ;
        RECT 1188.240000 371.420000 1189.980000 759.400000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1349.500000 2250.160000 1819.760000 2251.900000 ;
      LAYER met3 ;
        RECT 1349.500000 1863.920000 1819.760000 1865.660000 ;
      LAYER met4 ;
        RECT 1349.500000 1863.920000 1351.240000 2251.900000 ;
      LAYER met4 ;
        RECT 1818.020000 1863.920000 1819.760000 2251.900000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1349.500000 1752.660000 1819.760000 1754.400000 ;
      LAYER met3 ;
        RECT 1349.500000 1366.420000 1819.760000 1368.160000 ;
      LAYER met4 ;
        RECT 1349.500000 1366.420000 1351.240000 1754.400000 ;
      LAYER met4 ;
        RECT 1818.020000 1366.420000 1819.760000 1754.400000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1349.500000 1255.160000 1819.760000 1256.900000 ;
      LAYER met3 ;
        RECT 1349.500000 868.920000 1819.760000 870.660000 ;
      LAYER met4 ;
        RECT 1349.500000 868.920000 1351.240000 1256.900000 ;
      LAYER met4 ;
        RECT 1818.020000 868.920000 1819.760000 1256.900000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1349.500000 757.660000 1819.760000 759.400000 ;
      LAYER met3 ;
        RECT 1349.500000 371.420000 1819.760000 373.160000 ;
      LAYER met4 ;
        RECT 1349.500000 371.420000 1351.240000 759.400000 ;
      LAYER met4 ;
        RECT 1818.020000 371.420000 1819.760000 759.400000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1900.720000 2339.200000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1900.720000 2339.200000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 1900.720000 2339.200000 ;
    LAYER met3 ;
      RECT 1874.250000 2338.100000 1900.720000 2339.200000 ;
      RECT 1827.750000 2338.100000 1873.350000 2339.200000 ;
      RECT 1773.950000 2338.100000 1826.850000 2339.200000 ;
      RECT 1720.250000 2338.100000 1773.050000 2339.200000 ;
      RECT 1666.450000 2338.100000 1719.350000 2339.200000 ;
      RECT 1612.750000 2338.100000 1665.550000 2339.200000 ;
      RECT 1559.050000 2338.100000 1611.850000 2339.200000 ;
      RECT 1505.250000 2338.100000 1558.150000 2339.200000 ;
      RECT 1451.450000 2338.100000 1504.350000 2339.200000 ;
      RECT 1397.750000 2338.100000 1450.550000 2339.200000 ;
      RECT 1344.050000 2338.100000 1396.850000 2339.200000 ;
      RECT 1290.150000 2338.100000 1343.150000 2339.200000 ;
      RECT 1236.550000 2338.100000 1289.250000 2339.200000 ;
      RECT 1182.750000 2338.100000 1235.650000 2339.200000 ;
      RECT 1129.050000 2338.100000 1181.850000 2339.200000 ;
      RECT 1075.250000 2338.100000 1128.150000 2339.200000 ;
      RECT 1021.450000 2338.100000 1074.350000 2339.200000 ;
      RECT 967.850000 2338.100000 1020.550000 2339.200000 ;
      RECT 913.950000 2338.100000 966.950000 2339.200000 ;
      RECT 860.250000 2338.100000 913.050000 2339.200000 ;
      RECT 806.550000 2338.100000 859.350000 2339.200000 ;
      RECT 752.850000 2338.100000 805.650000 2339.200000 ;
      RECT 699.050000 2338.100000 751.950000 2339.200000 ;
      RECT 645.250000 2338.100000 698.150000 2339.200000 ;
      RECT 591.550000 2338.100000 644.350000 2339.200000 ;
      RECT 537.750000 2338.100000 590.650000 2339.200000 ;
      RECT 484.050000 2338.100000 536.850000 2339.200000 ;
      RECT 430.250000 2338.100000 483.150000 2339.200000 ;
      RECT 376.650000 2338.100000 429.350000 2339.200000 ;
      RECT 322.750000 2338.100000 375.750000 2339.200000 ;
      RECT 269.050000 2338.100000 321.850000 2339.200000 ;
      RECT 215.350000 2338.100000 268.150000 2339.200000 ;
      RECT 161.550000 2338.100000 214.450000 2339.200000 ;
      RECT 107.850000 2338.100000 160.650000 2339.200000 ;
      RECT 54.050000 2338.100000 106.950000 2339.200000 ;
      RECT 6.450000 2338.100000 53.150000 2339.200000 ;
      RECT 0.000000 2338.100000 5.550000 2339.200000 ;
      RECT 0.000000 1.100000 1900.720000 2338.100000 ;
      RECT 1878.850000 0.000000 1900.720000 1.100000 ;
      RECT 1876.150000 0.000000 1877.950000 1.100000 ;
      RECT 1873.450000 0.000000 1875.250000 1.100000 ;
      RECT 1869.650000 0.000000 1872.550000 1.100000 ;
      RECT 1865.950000 0.000000 1868.750000 1.100000 ;
      RECT 1862.050000 0.000000 1865.050000 1.100000 ;
      RECT 1858.150000 0.000000 1861.150000 1.100000 ;
      RECT 1854.450000 0.000000 1857.250000 1.100000 ;
      RECT 1850.650000 0.000000 1853.550000 1.100000 ;
      RECT 1846.850000 0.000000 1849.750000 1.100000 ;
      RECT 1842.950000 0.000000 1845.950000 1.100000 ;
      RECT 1839.150000 0.000000 1842.050000 1.100000 ;
      RECT 1835.350000 0.000000 1838.250000 1.100000 ;
      RECT 1831.550000 0.000000 1834.450000 1.100000 ;
      RECT 1827.750000 0.000000 1830.650000 1.100000 ;
      RECT 1823.850000 0.000000 1826.850000 1.100000 ;
      RECT 1820.050000 0.000000 1822.950000 1.100000 ;
      RECT 1816.350000 0.000000 1819.150000 1.100000 ;
      RECT 1812.450000 0.000000 1815.450000 1.100000 ;
      RECT 1808.550000 0.000000 1811.550000 1.100000 ;
      RECT 1804.850000 0.000000 1807.650000 1.100000 ;
      RECT 1801.050000 0.000000 1803.950000 1.100000 ;
      RECT 1797.250000 0.000000 1800.150000 1.100000 ;
      RECT 1793.350000 0.000000 1796.350000 1.100000 ;
      RECT 1789.550000 0.000000 1792.450000 1.100000 ;
      RECT 1785.750000 0.000000 1788.650000 1.100000 ;
      RECT 1781.950000 0.000000 1784.850000 1.100000 ;
      RECT 1778.050000 0.000000 1781.050000 1.100000 ;
      RECT 1774.350000 0.000000 1777.150000 1.100000 ;
      RECT 1770.450000 0.000000 1773.450000 1.100000 ;
      RECT 1766.750000 0.000000 1769.550000 1.100000 ;
      RECT 1762.850000 0.000000 1765.850000 1.100000 ;
      RECT 1759.050000 0.000000 1761.950000 1.100000 ;
      RECT 1755.250000 0.000000 1758.150000 1.100000 ;
      RECT 1751.450000 0.000000 1754.350000 1.100000 ;
      RECT 1747.550000 0.000000 1750.550000 1.100000 ;
      RECT 1743.750000 0.000000 1746.650000 1.100000 ;
      RECT 1739.950000 0.000000 1742.850000 1.100000 ;
      RECT 1736.150000 0.000000 1739.050000 1.100000 ;
      RECT 1732.350000 0.000000 1735.250000 1.100000 ;
      RECT 1728.450000 0.000000 1731.450000 1.100000 ;
      RECT 1724.750000 0.000000 1727.550000 1.100000 ;
      RECT 1720.850000 0.000000 1723.850000 1.100000 ;
      RECT 1717.150000 0.000000 1719.950000 1.100000 ;
      RECT 1713.250000 0.000000 1716.250000 1.100000 ;
      RECT 1709.450000 0.000000 1712.350000 1.100000 ;
      RECT 1705.650000 0.000000 1708.550000 1.100000 ;
      RECT 1701.850000 0.000000 1704.750000 1.100000 ;
      RECT 1697.950000 0.000000 1700.950000 1.100000 ;
      RECT 1694.250000 0.000000 1697.050000 1.100000 ;
      RECT 1690.350000 0.000000 1693.350000 1.100000 ;
      RECT 1686.550000 0.000000 1689.450000 1.100000 ;
      RECT 1682.750000 0.000000 1685.650000 1.100000 ;
      RECT 1678.950000 0.000000 1681.850000 1.100000 ;
      RECT 1675.150000 0.000000 1678.050000 1.100000 ;
      RECT 1671.250000 0.000000 1674.250000 1.100000 ;
      RECT 1667.450000 0.000000 1670.350000 1.100000 ;
      RECT 1663.650000 0.000000 1666.550000 1.100000 ;
      RECT 1659.850000 0.000000 1662.750000 1.100000 ;
      RECT 1656.050000 0.000000 1658.950000 1.100000 ;
      RECT 1652.250000 0.000000 1655.150000 1.100000 ;
      RECT 1648.350000 0.000000 1651.350000 1.100000 ;
      RECT 1644.650000 0.000000 1647.450000 1.100000 ;
      RECT 1640.750000 0.000000 1643.750000 1.100000 ;
      RECT 1636.950000 0.000000 1639.850000 1.100000 ;
      RECT 1633.150000 0.000000 1636.050000 1.100000 ;
      RECT 1629.350000 0.000000 1632.250000 1.100000 ;
      RECT 1625.550000 0.000000 1628.450000 1.100000 ;
      RECT 1621.650000 0.000000 1624.650000 1.100000 ;
      RECT 1617.850000 0.000000 1620.750000 1.100000 ;
      RECT 1614.150000 0.000000 1616.950000 1.100000 ;
      RECT 1610.250000 0.000000 1613.250000 1.100000 ;
      RECT 1606.450000 0.000000 1609.350000 1.100000 ;
      RECT 1602.650000 0.000000 1605.550000 1.100000 ;
      RECT 1598.850000 0.000000 1601.750000 1.100000 ;
      RECT 1595.050000 0.000000 1597.950000 1.100000 ;
      RECT 1591.150000 0.000000 1594.150000 1.100000 ;
      RECT 1587.250000 0.000000 1590.250000 1.100000 ;
      RECT 1583.550000 0.000000 1586.350000 1.100000 ;
      RECT 1579.750000 0.000000 1582.650000 1.100000 ;
      RECT 1575.950000 0.000000 1578.850000 1.100000 ;
      RECT 1572.050000 0.000000 1575.050000 1.100000 ;
      RECT 1568.250000 0.000000 1571.150000 1.100000 ;
      RECT 1564.550000 0.000000 1567.350000 1.100000 ;
      RECT 1560.650000 0.000000 1563.650000 1.100000 ;
      RECT 1556.750000 0.000000 1559.750000 1.100000 ;
      RECT 1553.050000 0.000000 1555.850000 1.100000 ;
      RECT 1549.250000 0.000000 1552.150000 1.100000 ;
      RECT 1545.450000 0.000000 1548.350000 1.100000 ;
      RECT 1541.550000 0.000000 1544.550000 1.100000 ;
      RECT 1537.650000 0.000000 1540.650000 1.100000 ;
      RECT 1534.050000 0.000000 1536.750000 1.100000 ;
      RECT 1530.150000 0.000000 1533.150000 1.100000 ;
      RECT 1526.350000 0.000000 1529.250000 1.100000 ;
      RECT 1522.450000 0.000000 1525.450000 1.100000 ;
      RECT 1518.750000 0.000000 1521.550000 1.100000 ;
      RECT 1514.950000 0.000000 1517.850000 1.100000 ;
      RECT 1511.050000 0.000000 1514.050000 1.100000 ;
      RECT 1507.150000 0.000000 1510.150000 1.100000 ;
      RECT 1503.450000 0.000000 1506.250000 1.100000 ;
      RECT 1499.650000 0.000000 1502.550000 1.100000 ;
      RECT 1495.850000 0.000000 1498.750000 1.100000 ;
      RECT 1491.950000 0.000000 1494.950000 1.100000 ;
      RECT 1488.150000 0.000000 1491.050000 1.100000 ;
      RECT 1484.450000 0.000000 1487.250000 1.100000 ;
      RECT 1480.550000 0.000000 1483.550000 1.100000 ;
      RECT 1476.650000 0.000000 1479.650000 1.100000 ;
      RECT 1472.850000 0.000000 1475.750000 1.100000 ;
      RECT 1469.150000 0.000000 1471.950000 1.100000 ;
      RECT 1465.350000 0.000000 1468.250000 1.100000 ;
      RECT 1461.450000 0.000000 1464.450000 1.100000 ;
      RECT 1457.550000 0.000000 1460.550000 1.100000 ;
      RECT 1453.950000 0.000000 1456.650000 1.100000 ;
      RECT 1450.050000 0.000000 1453.050000 1.100000 ;
      RECT 1446.250000 0.000000 1449.150000 1.100000 ;
      RECT 1442.350000 0.000000 1445.350000 1.100000 ;
      RECT 1438.550000 0.000000 1441.450000 1.100000 ;
      RECT 1434.850000 0.000000 1437.650000 1.100000 ;
      RECT 1430.950000 0.000000 1433.950000 1.100000 ;
      RECT 1427.050000 0.000000 1430.050000 1.100000 ;
      RECT 1423.350000 0.000000 1426.150000 1.100000 ;
      RECT 1419.550000 0.000000 1422.450000 1.100000 ;
      RECT 1415.750000 0.000000 1418.650000 1.100000 ;
      RECT 1411.850000 0.000000 1414.850000 1.100000 ;
      RECT 1408.050000 0.000000 1410.950000 1.100000 ;
      RECT 1404.350000 0.000000 1407.150000 1.100000 ;
      RECT 1400.450000 0.000000 1403.450000 1.100000 ;
      RECT 1396.550000 0.000000 1399.550000 1.100000 ;
      RECT 1392.750000 0.000000 1395.650000 1.100000 ;
      RECT 1388.950000 0.000000 1391.850000 1.100000 ;
      RECT 1385.250000 0.000000 1388.050000 1.100000 ;
      RECT 1381.350000 0.000000 1384.350000 1.100000 ;
      RECT 1377.450000 0.000000 1380.450000 1.100000 ;
      RECT 1373.750000 0.000000 1376.550000 1.100000 ;
      RECT 1369.950000 0.000000 1372.850000 1.100000 ;
      RECT 1366.050000 0.000000 1369.050000 1.100000 ;
      RECT 1362.250000 0.000000 1365.150000 1.100000 ;
      RECT 1358.450000 0.000000 1361.350000 1.100000 ;
      RECT 1354.750000 0.000000 1357.550000 1.100000 ;
      RECT 1350.850000 0.000000 1353.850000 1.100000 ;
      RECT 1346.950000 0.000000 1349.950000 1.100000 ;
      RECT 1343.250000 0.000000 1346.050000 1.100000 ;
      RECT 1339.350000 0.000000 1342.350000 1.100000 ;
      RECT 1335.650000 0.000000 1338.450000 1.100000 ;
      RECT 1331.750000 0.000000 1334.750000 1.100000 ;
      RECT 1327.950000 0.000000 1330.850000 1.100000 ;
      RECT 1324.150000 0.000000 1327.050000 1.100000 ;
      RECT 1320.350000 0.000000 1323.250000 1.100000 ;
      RECT 1316.450000 0.000000 1319.450000 1.100000 ;
      RECT 1312.650000 0.000000 1315.550000 1.100000 ;
      RECT 1308.850000 0.000000 1311.750000 1.100000 ;
      RECT 1305.150000 0.000000 1307.950000 1.100000 ;
      RECT 1301.250000 0.000000 1304.250000 1.100000 ;
      RECT 1297.350000 0.000000 1300.350000 1.100000 ;
      RECT 1293.650000 0.000000 1296.450000 1.100000 ;
      RECT 1289.750000 0.000000 1292.750000 1.100000 ;
      RECT 1285.950000 0.000000 1288.850000 1.100000 ;
      RECT 1282.150000 0.000000 1285.050000 1.100000 ;
      RECT 1278.350000 0.000000 1281.250000 1.100000 ;
      RECT 1274.550000 0.000000 1277.450000 1.100000 ;
      RECT 1270.750000 0.000000 1273.650000 1.100000 ;
      RECT 1266.850000 0.000000 1269.850000 1.100000 ;
      RECT 1263.150000 0.000000 1265.950000 1.100000 ;
      RECT 1259.250000 0.000000 1262.250000 1.100000 ;
      RECT 1255.550000 0.000000 1258.350000 1.100000 ;
      RECT 1251.650000 0.000000 1254.650000 1.100000 ;
      RECT 1247.850000 0.000000 1250.750000 1.100000 ;
      RECT 1244.050000 0.000000 1246.950000 1.100000 ;
      RECT 1240.150000 0.000000 1243.150000 1.100000 ;
      RECT 1236.350000 0.000000 1239.250000 1.100000 ;
      RECT 1232.550000 0.000000 1235.450000 1.100000 ;
      RECT 1228.750000 0.000000 1231.650000 1.100000 ;
      RECT 1224.950000 0.000000 1227.850000 1.100000 ;
      RECT 1221.150000 0.000000 1224.050000 1.100000 ;
      RECT 1217.250000 0.000000 1220.250000 1.100000 ;
      RECT 1213.550000 0.000000 1216.350000 1.100000 ;
      RECT 1209.650000 0.000000 1212.650000 1.100000 ;
      RECT 1205.850000 0.000000 1208.750000 1.100000 ;
      RECT 1202.050000 0.000000 1204.950000 1.100000 ;
      RECT 1198.250000 0.000000 1201.150000 1.100000 ;
      RECT 1194.450000 0.000000 1197.350000 1.100000 ;
      RECT 1190.550000 0.000000 1193.550000 1.100000 ;
      RECT 1186.750000 0.000000 1189.650000 1.100000 ;
      RECT 1183.050000 0.000000 1185.850000 1.100000 ;
      RECT 1179.150000 0.000000 1182.150000 1.100000 ;
      RECT 1175.250000 0.000000 1178.250000 1.100000 ;
      RECT 1171.550000 0.000000 1174.350000 1.100000 ;
      RECT 1167.750000 0.000000 1170.650000 1.100000 ;
      RECT 1163.950000 0.000000 1166.850000 1.100000 ;
      RECT 1160.050000 0.000000 1163.050000 1.100000 ;
      RECT 1156.250000 0.000000 1159.150000 1.100000 ;
      RECT 1152.450000 0.000000 1155.350000 1.100000 ;
      RECT 1148.650000 0.000000 1151.550000 1.100000 ;
      RECT 1144.850000 0.000000 1147.750000 1.100000 ;
      RECT 1140.950000 0.000000 1143.950000 1.100000 ;
      RECT 1137.150000 0.000000 1140.050000 1.100000 ;
      RECT 1133.450000 0.000000 1136.250000 1.100000 ;
      RECT 1129.550000 0.000000 1132.550000 1.100000 ;
      RECT 1125.650000 0.000000 1128.650000 1.100000 ;
      RECT 1121.950000 0.000000 1124.750000 1.100000 ;
      RECT 1118.150000 0.000000 1121.050000 1.100000 ;
      RECT 1114.350000 0.000000 1117.250000 1.100000 ;
      RECT 1110.450000 0.000000 1113.450000 1.100000 ;
      RECT 1106.650000 0.000000 1109.550000 1.100000 ;
      RECT 1102.950000 0.000000 1105.750000 1.100000 ;
      RECT 1099.050000 0.000000 1102.050000 1.100000 ;
      RECT 1095.150000 0.000000 1098.150000 1.100000 ;
      RECT 1091.350000 0.000000 1094.250000 1.100000 ;
      RECT 1087.650000 0.000000 1090.450000 1.100000 ;
      RECT 1083.850000 0.000000 1086.750000 1.100000 ;
      RECT 1079.950000 0.000000 1082.950000 1.100000 ;
      RECT 1076.050000 0.000000 1079.050000 1.100000 ;
      RECT 1072.350000 0.000000 1075.150000 1.100000 ;
      RECT 1068.550000 0.000000 1071.450000 1.100000 ;
      RECT 1064.750000 0.000000 1067.650000 1.100000 ;
      RECT 1060.850000 0.000000 1063.850000 1.100000 ;
      RECT 1057.050000 0.000000 1059.950000 1.100000 ;
      RECT 1053.350000 0.000000 1056.150000 1.100000 ;
      RECT 1049.450000 0.000000 1052.450000 1.100000 ;
      RECT 1045.550000 0.000000 1048.550000 1.100000 ;
      RECT 1041.750000 0.000000 1044.650000 1.100000 ;
      RECT 1038.050000 0.000000 1040.850000 1.100000 ;
      RECT 1034.250000 0.000000 1037.150000 1.100000 ;
      RECT 1030.350000 0.000000 1033.350000 1.100000 ;
      RECT 1026.450000 0.000000 1029.450000 1.100000 ;
      RECT 1022.850000 0.000000 1025.550000 1.100000 ;
      RECT 1018.950000 0.000000 1021.950000 1.100000 ;
      RECT 1015.050000 0.000000 1018.050000 1.100000 ;
      RECT 1011.250000 0.000000 1014.150000 1.100000 ;
      RECT 1007.550000 0.000000 1010.350000 1.100000 ;
      RECT 1003.750000 0.000000 1006.650000 1.100000 ;
      RECT 999.850000 0.000000 1002.850000 1.100000 ;
      RECT 995.950000 0.000000 998.950000 1.100000 ;
      RECT 992.250000 0.000000 995.050000 1.100000 ;
      RECT 988.450000 0.000000 991.350000 1.100000 ;
      RECT 984.550000 0.000000 987.550000 1.100000 ;
      RECT 980.750000 0.000000 983.650000 1.100000 ;
      RECT 976.950000 0.000000 979.850000 1.100000 ;
      RECT 973.250000 0.000000 976.050000 1.100000 ;
      RECT 969.350000 0.000000 972.350000 1.100000 ;
      RECT 965.450000 0.000000 968.450000 1.100000 ;
      RECT 961.650000 0.000000 964.550000 1.100000 ;
      RECT 957.950000 0.000000 960.750000 1.100000 ;
      RECT 954.150000 0.000000 957.050000 1.100000 ;
      RECT 950.250000 0.000000 953.250000 1.100000 ;
      RECT 946.350000 0.000000 949.350000 1.100000 ;
      RECT 942.650000 0.000000 945.450000 1.100000 ;
      RECT 938.850000 0.000000 941.750000 1.100000 ;
      RECT 934.950000 0.000000 937.950000 1.100000 ;
      RECT 931.150000 0.000000 934.050000 1.100000 ;
      RECT 927.350000 0.000000 930.250000 1.100000 ;
      RECT 923.650000 0.000000 926.450000 1.100000 ;
      RECT 919.750000 0.000000 922.750000 1.100000 ;
      RECT 915.850000 0.000000 918.850000 1.100000 ;
      RECT 912.150000 0.000000 914.950000 1.100000 ;
      RECT 908.350000 0.000000 911.250000 1.100000 ;
      RECT 904.450000 0.000000 907.450000 1.100000 ;
      RECT 900.650000 0.000000 903.550000 1.100000 ;
      RECT 896.850000 0.000000 899.750000 1.100000 ;
      RECT 893.050000 0.000000 895.950000 1.100000 ;
      RECT 889.250000 0.000000 892.150000 1.100000 ;
      RECT 885.350000 0.000000 888.350000 1.100000 ;
      RECT 881.550000 0.000000 884.450000 1.100000 ;
      RECT 877.750000 0.000000 880.650000 1.100000 ;
      RECT 874.050000 0.000000 876.850000 1.100000 ;
      RECT 870.150000 0.000000 873.150000 1.100000 ;
      RECT 866.250000 0.000000 869.250000 1.100000 ;
      RECT 862.550000 0.000000 865.350000 1.100000 ;
      RECT 858.750000 0.000000 861.650000 1.100000 ;
      RECT 854.850000 0.000000 857.850000 1.100000 ;
      RECT 851.050000 0.000000 853.950000 1.100000 ;
      RECT 847.250000 0.000000 850.150000 1.100000 ;
      RECT 843.450000 0.000000 846.350000 1.100000 ;
      RECT 839.650000 0.000000 842.550000 1.100000 ;
      RECT 835.750000 0.000000 838.750000 1.100000 ;
      RECT 832.050000 0.000000 834.850000 1.100000 ;
      RECT 828.150000 0.000000 831.150000 1.100000 ;
      RECT 824.350000 0.000000 827.250000 1.100000 ;
      RECT 820.550000 0.000000 823.450000 1.100000 ;
      RECT 816.750000 0.000000 819.650000 1.100000 ;
      RECT 812.950000 0.000000 815.850000 1.100000 ;
      RECT 809.150000 0.000000 812.050000 1.100000 ;
      RECT 805.250000 0.000000 808.250000 1.100000 ;
      RECT 801.450000 0.000000 804.350000 1.100000 ;
      RECT 797.650000 0.000000 800.550000 1.100000 ;
      RECT 793.850000 0.000000 796.750000 1.100000 ;
      RECT 790.050000 0.000000 792.950000 1.100000 ;
      RECT 786.150000 0.000000 789.150000 1.100000 ;
      RECT 782.450000 0.000000 785.250000 1.100000 ;
      RECT 778.550000 0.000000 781.550000 1.100000 ;
      RECT 774.750000 0.000000 777.650000 1.100000 ;
      RECT 770.950000 0.000000 773.850000 1.100000 ;
      RECT 767.150000 0.000000 770.050000 1.100000 ;
      RECT 763.350000 0.000000 766.250000 1.100000 ;
      RECT 759.550000 0.000000 762.450000 1.100000 ;
      RECT 755.650000 0.000000 758.650000 1.100000 ;
      RECT 751.950000 0.000000 754.750000 1.100000 ;
      RECT 748.050000 0.000000 751.050000 1.100000 ;
      RECT 744.250000 0.000000 747.150000 1.100000 ;
      RECT 740.450000 0.000000 743.350000 1.100000 ;
      RECT 736.650000 0.000000 739.550000 1.100000 ;
      RECT 732.850000 0.000000 735.750000 1.100000 ;
      RECT 728.950000 0.000000 731.950000 1.100000 ;
      RECT 725.150000 0.000000 728.050000 1.100000 ;
      RECT 721.350000 0.000000 724.250000 1.100000 ;
      RECT 717.550000 0.000000 720.450000 1.100000 ;
      RECT 713.650000 0.000000 716.650000 1.100000 ;
      RECT 709.950000 0.000000 712.750000 1.100000 ;
      RECT 706.050000 0.000000 709.050000 1.100000 ;
      RECT 702.350000 0.000000 705.150000 1.100000 ;
      RECT 698.450000 0.000000 701.450000 1.100000 ;
      RECT 694.650000 0.000000 697.550000 1.100000 ;
      RECT 690.850000 0.000000 693.750000 1.100000 ;
      RECT 687.050000 0.000000 689.950000 1.100000 ;
      RECT 683.250000 0.000000 686.150000 1.100000 ;
      RECT 679.350000 0.000000 682.350000 1.100000 ;
      RECT 675.550000 0.000000 678.450000 1.100000 ;
      RECT 671.850000 0.000000 674.650000 1.100000 ;
      RECT 667.950000 0.000000 670.950000 1.100000 ;
      RECT 664.050000 0.000000 667.050000 1.100000 ;
      RECT 660.350000 0.000000 663.150000 1.100000 ;
      RECT 656.550000 0.000000 659.450000 1.100000 ;
      RECT 652.750000 0.000000 655.650000 1.100000 ;
      RECT 648.850000 0.000000 651.850000 1.100000 ;
      RECT 645.050000 0.000000 647.950000 1.100000 ;
      RECT 641.250000 0.000000 644.150000 1.100000 ;
      RECT 637.450000 0.000000 640.350000 1.100000 ;
      RECT 633.550000 0.000000 636.550000 1.100000 ;
      RECT 629.750000 0.000000 632.650000 1.100000 ;
      RECT 625.950000 0.000000 628.850000 1.100000 ;
      RECT 622.250000 0.000000 625.050000 1.100000 ;
      RECT 618.350000 0.000000 621.350000 1.100000 ;
      RECT 614.450000 0.000000 617.450000 1.100000 ;
      RECT 610.750000 0.000000 613.550000 1.100000 ;
      RECT 606.950000 0.000000 609.850000 1.100000 ;
      RECT 603.050000 0.000000 606.050000 1.100000 ;
      RECT 599.250000 0.000000 602.150000 1.100000 ;
      RECT 595.450000 0.000000 598.350000 1.100000 ;
      RECT 591.750000 0.000000 594.550000 1.100000 ;
      RECT 587.850000 0.000000 590.850000 1.100000 ;
      RECT 583.950000 0.000000 586.950000 1.100000 ;
      RECT 580.150000 0.000000 583.050000 1.100000 ;
      RECT 576.450000 0.000000 579.250000 1.100000 ;
      RECT 572.650000 0.000000 575.550000 1.100000 ;
      RECT 568.750000 0.000000 571.750000 1.100000 ;
      RECT 564.850000 0.000000 567.850000 1.100000 ;
      RECT 561.150000 0.000000 563.950000 1.100000 ;
      RECT 557.350000 0.000000 560.250000 1.100000 ;
      RECT 553.450000 0.000000 556.450000 1.100000 ;
      RECT 549.650000 0.000000 552.550000 1.100000 ;
      RECT 545.850000 0.000000 548.750000 1.100000 ;
      RECT 542.150000 0.000000 544.950000 1.100000 ;
      RECT 538.250000 0.000000 541.250000 1.100000 ;
      RECT 534.350000 0.000000 537.350000 1.100000 ;
      RECT 530.550000 0.000000 533.450000 1.100000 ;
      RECT 526.850000 0.000000 529.650000 1.100000 ;
      RECT 522.950000 0.000000 525.950000 1.100000 ;
      RECT 519.150000 0.000000 522.050000 1.100000 ;
      RECT 515.250000 0.000000 518.250000 1.100000 ;
      RECT 511.650000 0.000000 514.350000 1.100000 ;
      RECT 507.750000 0.000000 510.750000 1.100000 ;
      RECT 503.850000 0.000000 506.850000 1.100000 ;
      RECT 500.050000 0.000000 502.950000 1.100000 ;
      RECT 496.350000 0.000000 499.150000 1.100000 ;
      RECT 492.550000 0.000000 495.450000 1.100000 ;
      RECT 488.650000 0.000000 491.650000 1.100000 ;
      RECT 484.750000 0.000000 487.750000 1.100000 ;
      RECT 481.050000 0.000000 483.850000 1.100000 ;
      RECT 477.250000 0.000000 480.150000 1.100000 ;
      RECT 473.350000 0.000000 476.350000 1.100000 ;
      RECT 469.550000 0.000000 472.450000 1.100000 ;
      RECT 465.750000 0.000000 468.650000 1.100000 ;
      RECT 462.050000 0.000000 464.850000 1.100000 ;
      RECT 458.150000 0.000000 461.150000 1.100000 ;
      RECT 454.250000 0.000000 457.250000 1.100000 ;
      RECT 450.450000 0.000000 453.350000 1.100000 ;
      RECT 446.750000 0.000000 449.550000 1.100000 ;
      RECT 442.850000 0.000000 445.850000 1.100000 ;
      RECT 439.050000 0.000000 441.950000 1.100000 ;
      RECT 435.150000 0.000000 438.150000 1.100000 ;
      RECT 431.450000 0.000000 434.250000 1.100000 ;
      RECT 427.650000 0.000000 430.550000 1.100000 ;
      RECT 423.750000 0.000000 426.750000 1.100000 ;
      RECT 419.950000 0.000000 422.850000 1.100000 ;
      RECT 416.150000 0.000000 419.050000 1.100000 ;
      RECT 412.350000 0.000000 415.250000 1.100000 ;
      RECT 408.550000 0.000000 411.450000 1.100000 ;
      RECT 404.650000 0.000000 407.650000 1.100000 ;
      RECT 400.950000 0.000000 403.750000 1.100000 ;
      RECT 397.150000 0.000000 400.050000 1.100000 ;
      RECT 393.250000 0.000000 396.250000 1.100000 ;
      RECT 389.450000 0.000000 392.350000 1.100000 ;
      RECT 385.650000 0.000000 388.550000 1.100000 ;
      RECT 381.850000 0.000000 384.750000 1.100000 ;
      RECT 378.050000 0.000000 380.950000 1.100000 ;
      RECT 374.150000 0.000000 377.150000 1.100000 ;
      RECT 370.350000 0.000000 373.250000 1.100000 ;
      RECT 366.550000 0.000000 369.450000 1.100000 ;
      RECT 362.750000 0.000000 365.650000 1.100000 ;
      RECT 358.950000 0.000000 361.850000 1.100000 ;
      RECT 355.050000 0.000000 358.050000 1.100000 ;
      RECT 351.350000 0.000000 354.150000 1.100000 ;
      RECT 347.550000 0.000000 350.450000 1.100000 ;
      RECT 343.650000 0.000000 346.650000 1.100000 ;
      RECT 339.850000 0.000000 342.750000 1.100000 ;
      RECT 336.050000 0.000000 338.950000 1.100000 ;
      RECT 332.150000 0.000000 335.150000 1.100000 ;
      RECT 328.450000 0.000000 331.250000 1.100000 ;
      RECT 324.550000 0.000000 327.550000 1.100000 ;
      RECT 320.850000 0.000000 323.650000 1.100000 ;
      RECT 316.950000 0.000000 319.950000 1.100000 ;
      RECT 313.150000 0.000000 316.050000 1.100000 ;
      RECT 309.350000 0.000000 312.250000 1.100000 ;
      RECT 305.550000 0.000000 308.450000 1.100000 ;
      RECT 301.750000 0.000000 304.650000 1.100000 ;
      RECT 297.950000 0.000000 300.850000 1.100000 ;
      RECT 294.050000 0.000000 297.050000 1.100000 ;
      RECT 290.250000 0.000000 293.150000 1.100000 ;
      RECT 286.450000 0.000000 289.350000 1.100000 ;
      RECT 282.550000 0.000000 285.550000 1.100000 ;
      RECT 278.850000 0.000000 281.650000 1.100000 ;
      RECT 274.950000 0.000000 277.950000 1.100000 ;
      RECT 271.250000 0.000000 274.050000 1.100000 ;
      RECT 267.350000 0.000000 270.350000 1.100000 ;
      RECT 263.550000 0.000000 266.450000 1.100000 ;
      RECT 259.750000 0.000000 262.650000 1.100000 ;
      RECT 255.950000 0.000000 258.850000 1.100000 ;
      RECT 252.050000 0.000000 255.050000 1.100000 ;
      RECT 248.350000 0.000000 251.150000 1.100000 ;
      RECT 244.450000 0.000000 247.450000 1.100000 ;
      RECT 240.750000 0.000000 243.550000 1.100000 ;
      RECT 236.850000 0.000000 239.850000 1.100000 ;
      RECT 232.950000 0.000000 235.950000 1.100000 ;
      RECT 229.250000 0.000000 232.050000 1.100000 ;
      RECT 225.450000 0.000000 228.350000 1.100000 ;
      RECT 221.550000 0.000000 224.550000 1.100000 ;
      RECT 217.750000 0.000000 220.650000 1.100000 ;
      RECT 213.950000 0.000000 216.850000 1.100000 ;
      RECT 210.150000 0.000000 213.050000 1.100000 ;
      RECT 206.350000 0.000000 209.250000 1.100000 ;
      RECT 202.450000 0.000000 205.450000 1.100000 ;
      RECT 198.750000 0.000000 201.550000 1.100000 ;
      RECT 194.850000 0.000000 197.850000 1.100000 ;
      RECT 191.150000 0.000000 193.950000 1.100000 ;
      RECT 187.250000 0.000000 190.250000 1.100000 ;
      RECT 183.350000 0.000000 186.350000 1.100000 ;
      RECT 179.650000 0.000000 182.450000 1.100000 ;
      RECT 175.850000 0.000000 178.750000 1.100000 ;
      RECT 171.950000 0.000000 174.950000 1.100000 ;
      RECT 168.150000 0.000000 171.050000 1.100000 ;
      RECT 164.350000 0.000000 167.250000 1.100000 ;
      RECT 160.650000 0.000000 163.450000 1.100000 ;
      RECT 156.750000 0.000000 159.750000 1.100000 ;
      RECT 152.850000 0.000000 155.850000 1.100000 ;
      RECT 149.150000 0.000000 151.950000 1.100000 ;
      RECT 145.350000 0.000000 148.250000 1.100000 ;
      RECT 141.450000 0.000000 144.450000 1.100000 ;
      RECT 137.650000 0.000000 140.550000 1.100000 ;
      RECT 133.750000 0.000000 136.750000 1.100000 ;
      RECT 130.050000 0.000000 132.850000 1.100000 ;
      RECT 126.250000 0.000000 129.150000 1.100000 ;
      RECT 122.350000 0.000000 125.350000 1.100000 ;
      RECT 118.550000 0.000000 121.450000 1.100000 ;
      RECT 114.750000 0.000000 117.650000 1.100000 ;
      RECT 111.050000 0.000000 113.850000 1.100000 ;
      RECT 107.150000 0.000000 110.150000 1.100000 ;
      RECT 103.250000 0.000000 106.250000 1.100000 ;
      RECT 99.550000 0.000000 102.350000 1.100000 ;
      RECT 95.750000 0.000000 98.650000 1.100000 ;
      RECT 91.850000 0.000000 94.850000 1.100000 ;
      RECT 88.050000 0.000000 90.950000 1.100000 ;
      RECT 84.150000 0.000000 87.150000 1.100000 ;
      RECT 80.550000 0.000000 83.250000 1.100000 ;
      RECT 76.650000 0.000000 79.650000 1.100000 ;
      RECT 72.750000 0.000000 75.750000 1.100000 ;
      RECT 68.950000 0.000000 71.850000 1.100000 ;
      RECT 65.250000 0.000000 68.050000 1.100000 ;
      RECT 61.350000 0.000000 64.350000 1.100000 ;
      RECT 57.550000 0.000000 60.450000 1.100000 ;
      RECT 53.650000 0.000000 56.650000 1.100000 ;
      RECT 49.950000 0.000000 52.750000 1.100000 ;
      RECT 46.150000 0.000000 49.050000 1.100000 ;
      RECT 42.250000 0.000000 45.250000 1.100000 ;
      RECT 38.450000 0.000000 41.350000 1.100000 ;
      RECT 34.650000 0.000000 37.550000 1.100000 ;
      RECT 30.850000 0.000000 33.750000 1.100000 ;
      RECT 27.050000 0.000000 29.950000 1.100000 ;
      RECT 23.150000 0.000000 26.150000 1.100000 ;
      RECT 19.350000 0.000000 22.250000 1.100000 ;
      RECT 15.650000 0.000000 18.450000 1.100000 ;
      RECT 11.750000 0.000000 14.750000 1.100000 ;
      RECT 7.950000 0.000000 10.850000 1.100000 ;
      RECT 5.650000 0.000000 7.050000 1.100000 ;
      RECT 2.150000 0.000000 4.750000 1.100000 ;
      RECT 0.000000 0.000000 1.250000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 2330.860000 1900.720000 2339.200000 ;
      RECT 12.180000 2324.860000 1888.080000 2330.860000 ;
      RECT 1892.880000 2308.045000 1900.720000 2330.860000 ;
      RECT 0.000000 2307.125000 7.380000 2330.860000 ;
      RECT 1892.880000 2307.045000 1899.620000 2308.045000 ;
      RECT 1.100000 2306.125000 7.380000 2307.125000 ;
      RECT 0.000000 2270.140000 7.380000 2306.125000 ;
      RECT 1892.880000 2269.310000 1900.720000 2307.045000 ;
      RECT 1.100000 2269.140000 7.380000 2270.140000 ;
      RECT 1892.880000 2268.310000 1899.620000 2269.310000 ;
      RECT 0.000000 2226.530000 7.380000 2269.140000 ;
      RECT 1.100000 2225.530000 7.380000 2226.530000 ;
      RECT 1892.880000 2224.785000 1900.720000 2268.310000 ;
      RECT 1892.880000 2223.785000 1899.620000 2224.785000 ;
      RECT 0.000000 2182.925000 7.380000 2225.530000 ;
      RECT 1.100000 2181.925000 7.380000 2182.925000 ;
      RECT 1892.880000 2180.255000 1900.720000 2223.785000 ;
      RECT 1892.880000 2179.255000 1899.620000 2180.255000 ;
      RECT 0.000000 2139.225000 7.380000 2181.925000 ;
      RECT 1.100000 2138.225000 7.380000 2139.225000 ;
      RECT 1892.880000 2135.820000 1900.720000 2179.255000 ;
      RECT 1892.880000 2134.820000 1899.620000 2135.820000 ;
      RECT 0.000000 2095.430000 7.380000 2138.225000 ;
      RECT 1.100000 2094.430000 7.380000 2095.430000 ;
      RECT 1892.880000 2091.290000 1900.720000 2134.820000 ;
      RECT 1892.880000 2090.290000 1899.620000 2091.290000 ;
      RECT 0.000000 2051.915000 7.380000 2094.430000 ;
      RECT 1.100000 2050.915000 7.380000 2051.915000 ;
      RECT 1892.880000 2046.855000 1900.720000 2090.290000 ;
      RECT 1892.880000 2045.855000 1899.620000 2046.855000 ;
      RECT 0.000000 2008.215000 7.380000 2050.915000 ;
      RECT 1.100000 2007.215000 7.380000 2008.215000 ;
      RECT 1892.880000 2002.330000 1900.720000 2045.855000 ;
      RECT 1892.880000 2001.330000 1899.620000 2002.330000 ;
      RECT 0.000000 1964.610000 7.380000 2007.215000 ;
      RECT 1.100000 1963.610000 7.380000 1964.610000 ;
      RECT 1892.880000 1957.800000 1900.720000 2001.330000 ;
      RECT 1892.880000 1956.800000 1899.620000 1957.800000 ;
      RECT 0.000000 1920.910000 7.380000 1963.610000 ;
      RECT 1.100000 1919.910000 7.380000 1920.910000 ;
      RECT 1892.880000 1913.365000 1900.720000 1956.800000 ;
      RECT 1892.880000 1912.365000 1899.620000 1913.365000 ;
      RECT 0.000000 1877.300000 7.380000 1919.910000 ;
      RECT 1.100000 1876.300000 7.380000 1877.300000 ;
      RECT 1892.880000 1868.930000 1900.720000 1912.365000 ;
      RECT 1892.880000 1867.930000 1899.620000 1868.930000 ;
      RECT 0.000000 1833.600000 7.380000 1876.300000 ;
      RECT 1.100000 1832.600000 7.380000 1833.600000 ;
      RECT 1892.880000 1824.400000 1900.720000 1867.930000 ;
      RECT 1892.880000 1823.400000 1899.620000 1824.400000 ;
      RECT 0.000000 1789.990000 7.380000 1832.600000 ;
      RECT 1.100000 1788.990000 7.380000 1789.990000 ;
      RECT 1892.880000 1779.965000 1900.720000 1823.400000 ;
      RECT 1892.880000 1778.965000 1899.620000 1779.965000 ;
      RECT 0.000000 1746.290000 7.380000 1788.990000 ;
      RECT 1.100000 1745.290000 7.380000 1746.290000 ;
      RECT 1892.880000 1735.530000 1900.720000 1778.965000 ;
      RECT 1892.880000 1734.530000 1899.620000 1735.530000 ;
      RECT 0.000000 1702.775000 7.380000 1745.290000 ;
      RECT 1.100000 1701.775000 7.380000 1702.775000 ;
      RECT 1892.880000 1690.910000 1900.720000 1734.530000 ;
      RECT 1892.880000 1689.910000 1899.620000 1690.910000 ;
      RECT 0.000000 1659.075000 7.380000 1701.775000 ;
      RECT 1.100000 1658.075000 7.380000 1659.075000 ;
      RECT 1892.880000 1646.470000 1900.720000 1689.910000 ;
      RECT 1892.880000 1645.470000 1899.620000 1646.470000 ;
      RECT 0.000000 1615.375000 7.380000 1658.075000 ;
      RECT 1.100000 1614.375000 7.380000 1615.375000 ;
      RECT 1892.880000 1601.945000 1900.720000 1645.470000 ;
      RECT 1892.880000 1600.945000 1899.620000 1601.945000 ;
      RECT 0.000000 1571.675000 7.380000 1614.375000 ;
      RECT 1.100000 1570.675000 7.380000 1571.675000 ;
      RECT 1892.880000 1557.510000 1900.720000 1600.945000 ;
      RECT 1892.880000 1556.510000 1899.620000 1557.510000 ;
      RECT 0.000000 1528.160000 7.380000 1570.675000 ;
      RECT 1.100000 1527.160000 7.380000 1528.160000 ;
      RECT 1892.880000 1512.980000 1900.720000 1556.510000 ;
      RECT 1892.880000 1511.980000 1899.620000 1512.980000 ;
      RECT 0.000000 1484.460000 7.380000 1527.160000 ;
      RECT 1.100000 1483.460000 7.380000 1484.460000 ;
      RECT 1892.880000 1468.450000 1900.720000 1511.980000 ;
      RECT 1892.880000 1467.450000 1899.620000 1468.450000 ;
      RECT 0.000000 1440.850000 7.380000 1483.460000 ;
      RECT 1.100000 1439.850000 7.380000 1440.850000 ;
      RECT 1892.880000 1424.015000 1900.720000 1467.450000 ;
      RECT 1892.880000 1423.015000 1899.620000 1424.015000 ;
      RECT 0.000000 1397.060000 7.380000 1439.850000 ;
      RECT 1.100000 1396.060000 7.380000 1397.060000 ;
      RECT 1892.880000 1379.490000 1900.720000 1423.015000 ;
      RECT 1892.880000 1378.490000 1899.620000 1379.490000 ;
      RECT 0.000000 1353.545000 7.380000 1396.060000 ;
      RECT 1.100000 1352.545000 7.380000 1353.545000 ;
      RECT 1892.880000 1335.050000 1900.720000 1378.490000 ;
      RECT 1892.880000 1334.050000 1899.620000 1335.050000 ;
      RECT 0.000000 1309.845000 7.380000 1352.545000 ;
      RECT 1.100000 1308.845000 7.380000 1309.845000 ;
      RECT 1892.880000 1290.525000 1900.720000 1334.050000 ;
      RECT 1892.880000 1289.525000 1899.620000 1290.525000 ;
      RECT 0.000000 1266.235000 7.380000 1308.845000 ;
      RECT 1.100000 1265.235000 7.380000 1266.235000 ;
      RECT 1892.880000 1246.090000 1900.720000 1289.525000 ;
      RECT 1892.880000 1245.090000 1899.620000 1246.090000 ;
      RECT 0.000000 1222.535000 7.380000 1265.235000 ;
      RECT 1.100000 1221.535000 7.380000 1222.535000 ;
      RECT 1892.880000 1201.470000 1900.720000 1245.090000 ;
      RECT 1892.880000 1200.470000 1899.620000 1201.470000 ;
      RECT 0.000000 1178.930000 7.380000 1221.535000 ;
      RECT 1.100000 1177.930000 7.380000 1178.930000 ;
      RECT 1892.880000 1157.030000 1900.720000 1200.470000 ;
      RECT 1892.880000 1156.030000 1899.620000 1157.030000 ;
      RECT 0.000000 1135.230000 7.380000 1177.930000 ;
      RECT 1.100000 1134.230000 7.380000 1135.230000 ;
      RECT 1892.880000 1112.505000 1900.720000 1156.030000 ;
      RECT 1892.880000 1111.505000 1899.620000 1112.505000 ;
      RECT 0.000000 1091.620000 7.380000 1134.230000 ;
      RECT 1.100000 1090.620000 7.380000 1091.620000 ;
      RECT 1892.880000 1068.070000 1900.720000 1111.505000 ;
      RECT 1892.880000 1067.070000 1899.620000 1068.070000 ;
      RECT 0.000000 1047.920000 7.380000 1090.620000 ;
      RECT 1.100000 1046.920000 7.380000 1047.920000 ;
      RECT 1892.880000 1023.630000 1900.720000 1067.070000 ;
      RECT 1892.880000 1022.630000 1899.620000 1023.630000 ;
      RECT 0.000000 1004.310000 7.380000 1046.920000 ;
      RECT 1.100000 1003.310000 7.380000 1004.310000 ;
      RECT 1892.880000 979.105000 1900.720000 1022.630000 ;
      RECT 1892.880000 978.105000 1899.620000 979.105000 ;
      RECT 0.000000 960.705000 7.380000 1003.310000 ;
      RECT 1.100000 959.705000 7.380000 960.705000 ;
      RECT 1892.880000 934.670000 1900.720000 978.105000 ;
      RECT 1892.880000 933.670000 1899.620000 934.670000 ;
      RECT 0.000000 916.910000 7.380000 959.705000 ;
      RECT 1.100000 915.910000 7.380000 916.910000 ;
      RECT 1892.880000 890.140000 1900.720000 933.670000 ;
      RECT 1892.880000 889.140000 1899.620000 890.140000 ;
      RECT 0.000000 873.305000 7.380000 915.910000 ;
      RECT 1.100000 872.305000 7.380000 873.305000 ;
      RECT 1892.880000 845.705000 1900.720000 889.140000 ;
      RECT 1892.880000 844.705000 1899.620000 845.705000 ;
      RECT 0.000000 829.695000 7.380000 872.305000 ;
      RECT 1.100000 828.695000 7.380000 829.695000 ;
      RECT 1892.880000 801.175000 1900.720000 844.705000 ;
      RECT 1892.880000 800.175000 1899.620000 801.175000 ;
      RECT 0.000000 786.090000 7.380000 828.695000 ;
      RECT 1.100000 785.090000 7.380000 786.090000 ;
      RECT 1892.880000 756.740000 1900.720000 800.175000 ;
      RECT 1892.880000 755.740000 1899.620000 756.740000 ;
      RECT 0.000000 742.390000 7.380000 785.090000 ;
      RECT 1.100000 741.390000 7.380000 742.390000 ;
      RECT 1892.880000 712.210000 1900.720000 755.740000 ;
      RECT 1892.880000 711.210000 1899.620000 712.210000 ;
      RECT 0.000000 698.780000 7.380000 741.390000 ;
      RECT 1.100000 697.780000 7.380000 698.780000 ;
      RECT 1892.880000 667.685000 1900.720000 711.210000 ;
      RECT 1892.880000 666.685000 1899.620000 667.685000 ;
      RECT 0.000000 655.080000 7.380000 697.780000 ;
      RECT 1.100000 654.080000 7.380000 655.080000 ;
      RECT 1892.880000 623.250000 1900.720000 666.685000 ;
      RECT 1892.880000 622.250000 1899.620000 623.250000 ;
      RECT 0.000000 611.470000 7.380000 654.080000 ;
      RECT 1.100000 610.470000 7.380000 611.470000 ;
      RECT 1892.880000 578.720000 1900.720000 622.250000 ;
      RECT 1892.880000 577.720000 1899.620000 578.720000 ;
      RECT 0.000000 567.770000 7.380000 610.470000 ;
      RECT 1.100000 566.770000 7.380000 567.770000 ;
      RECT 1892.880000 534.285000 1900.720000 577.720000 ;
      RECT 1892.880000 533.285000 1899.620000 534.285000 ;
      RECT 0.000000 524.165000 7.380000 566.770000 ;
      RECT 1.100000 523.165000 7.380000 524.165000 ;
      RECT 1892.880000 489.755000 1900.720000 533.285000 ;
      RECT 1892.880000 488.755000 1899.620000 489.755000 ;
      RECT 0.000000 480.555000 7.380000 523.165000 ;
      RECT 1.100000 479.555000 7.380000 480.555000 ;
      RECT 1892.880000 445.230000 1900.720000 488.755000 ;
      RECT 1892.880000 444.230000 1899.620000 445.230000 ;
      RECT 0.000000 436.855000 7.380000 479.555000 ;
      RECT 1.100000 435.855000 7.380000 436.855000 ;
      RECT 1892.880000 400.790000 1900.720000 444.230000 ;
      RECT 1892.880000 399.790000 1899.620000 400.790000 ;
      RECT 0.000000 393.155000 7.380000 435.855000 ;
      RECT 1.100000 392.155000 7.380000 393.155000 ;
      RECT 1892.880000 356.265000 1900.720000 399.790000 ;
      RECT 1892.880000 355.265000 1899.620000 356.265000 ;
      RECT 0.000000 349.640000 7.380000 392.155000 ;
      RECT 1.100000 348.640000 7.380000 349.640000 ;
      RECT 1892.880000 311.830000 1900.720000 355.265000 ;
      RECT 1892.880000 310.830000 1899.620000 311.830000 ;
      RECT 0.000000 305.940000 7.380000 348.640000 ;
      RECT 1.100000 304.940000 7.380000 305.940000 ;
      RECT 1892.880000 267.300000 1900.720000 310.830000 ;
      RECT 1892.880000 266.300000 1899.620000 267.300000 ;
      RECT 0.000000 262.330000 7.380000 304.940000 ;
      RECT 1.100000 261.330000 7.380000 262.330000 ;
      RECT 1892.880000 222.770000 1900.720000 266.300000 ;
      RECT 1892.880000 221.770000 1899.620000 222.770000 ;
      RECT 0.000000 218.540000 7.380000 261.330000 ;
      RECT 1.100000 217.540000 7.380000 218.540000 ;
      RECT 1892.880000 178.245000 1900.720000 221.770000 ;
      RECT 1892.880000 177.245000 1899.620000 178.245000 ;
      RECT 0.000000 175.025000 7.380000 217.540000 ;
      RECT 1.100000 174.025000 7.380000 175.025000 ;
      RECT 1892.880000 133.810000 1900.720000 177.245000 ;
      RECT 1892.880000 132.810000 1899.620000 133.810000 ;
      RECT 0.000000 131.325000 7.380000 174.025000 ;
      RECT 1.100000 130.325000 7.380000 131.325000 ;
      RECT 1892.880000 89.370000 1900.720000 132.810000 ;
      RECT 1892.880000 88.370000 1899.620000 89.370000 ;
      RECT 0.000000 87.715000 7.380000 130.325000 ;
      RECT 1.100000 86.715000 7.380000 87.715000 ;
      RECT 1892.880000 44.935000 1900.720000 88.370000 ;
      RECT 0.000000 44.015000 7.380000 86.715000 ;
      RECT 1892.880000 43.935000 1899.620000 44.935000 ;
      RECT 1.100000 43.015000 7.380000 44.015000 ;
      RECT 1886.880000 13.660000 1888.080000 2324.860000 ;
      RECT 18.180000 13.660000 1882.080000 2324.860000 ;
      RECT 12.180000 13.660000 13.380000 2324.860000 ;
      RECT 1892.880000 11.540000 1900.720000 43.935000 ;
      RECT 1892.880000 10.540000 1899.620000 11.540000 ;
      RECT 1892.880000 7.660000 1900.720000 10.540000 ;
      RECT 12.180000 7.660000 1888.080000 13.660000 ;
      RECT 0.000000 7.660000 7.380000 43.015000 ;
      RECT 0.000000 4.730000 1900.720000 7.660000 ;
      RECT 1.100000 3.730000 1900.720000 4.730000 ;
      RECT 0.000000 0.000000 1900.720000 3.730000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
